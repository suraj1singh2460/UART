library verilog;
use verilog.vl_types.all;
entity uart_pkg is
end uart_pkg;
