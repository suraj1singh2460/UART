library verilog;
use verilog.vl_types.all;
entity param_pkg is
end param_pkg;
